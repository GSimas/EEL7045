** Profile: "SCHEMATIC1-NewSim"  [ C:\USERS\GUSTAVO\DOCUMENTS\UFSC\4� FASE\CIRCUITOS EL�TRICOS A\EEL7045\Simulacoes\exemplo-SCHEMATIC1-NewSim.sim ] 

** Creating circuit file "exemplo-SCHEMATIC1-NewSim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 
.PROBE 
.INC "exemplo-SCHEMATIC1.net" 

.INC "exemplo-SCHEMATIC1.als"


.END
