** Profile: "SCHEMATIC1-NewSim"  [ C:\USERS\GUSTAVO\DOCUMENTS\UFSC\4� FASE\CIRCUITOS EL�TRICOS A\EEL7045\Simulacoes\rlc_serie-SCHEMATIC1-NewSim.sim ] 

** Creating circuit file "rlc_serie-SCHEMATIC1-NewSim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 4s 0 
.PROBE 
.INC "rlc_serie-SCHEMATIC1.net" 

.INC "rlc_serie-SCHEMATIC1.als"


.END
